`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:30:38 03/19/2020 
// Design Name: 
// Module Name:    microcode_executor 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module microcode_executor(
    input [7:0] r_addr,
    input [7:0] w_addr,
    inout [7:0] bus,
    input clk
    );


endmodule
