`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:28:55 03/19/2020 
// Design Name: 
// Module Name:    io_mem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module io_mem(
    input [7:0] r_addr,
    input [7:0] w_addr,
    inout [7:0] bus,
    input clk
    );


endmodule
